`timescale 1ns / 1ps

module ins_storage(
     address,dataout
    );
    input [11:0]address;
    output reg [31:0]dataout;
    reg [31:0]data[0:4095];
    initial 
    begin
    data[0]=32'h20110001;
    data[1]=32'h08000005;
    data[2]=32'h20110001;
    data[3]=32'h20120002;
    data[4]=32'h20130003;
    data[5]=32'h08000c09;
    data[6]=32'h20110001;
    data[7]=32'h20120002;
    data[8]=32'h20130003;
    data[9]=32'h0800000d;
    data[10]=32'h20110001;
    data[11]=32'h20120002;
    data[12]=32'h20130003;
    data[13]=32'h08000011;
    data[14]=32'h20110001;
    data[15]=32'h20120002;
    data[16]=32'h20130003;
    data[17]=32'h0c0000b8;
    data[18]=32'h20100001;
    data[19]=32'h20110001;
    data[20]=32'h00118fc0;
    data[21]=32'h00112020;
    data[22]=32'h20020022;
    data[23]=32'h0000000c;
    data[24]=32'h00118882;
    data[25]=32'h12200001;
    data[26]=32'h08000015;
    data[27]=32'h00112020;
    data[28]=32'h20020022;
    data[29]=32'h0000000c;
    data[30]=32'h20110001;
    data[31]=32'h00118880;
    data[32]=32'h00112020;
    data[33]=32'h20020022;
    data[34]=32'h0000000c;
    data[35]=32'h12200001;
    data[36]=32'h0800001f;
    data[37]=32'h20110001;
    data[38]=32'h00118fc0;
    data[39]=32'h00112020;
    data[40]=32'h20020022;
    data[41]=32'h0000000c;
    data[42]=32'h001188c3;
    data[43]=32'h00112020;
    data[44]=32'h20020022;
    data[45]=32'h0000000c;
    data[46]=32'h00118903;
    data[47]=32'h00112020;
    data[48]=32'h20020022;
    data[49]=32'h0000000c;
    data[50]=32'h00118903;
    data[51]=32'h00112020;
    data[52]=32'h20020022;
    data[53]=32'h0000000c;
    data[54]=32'h00118903;
    data[55]=32'h00112020;
    data[56]=32'h20020022;
    data[57]=32'h0000000c;
    data[58]=32'h00118903;
    data[59]=32'h00112020;
    data[60]=32'h20020022;
    data[61]=32'h0000000c;
    data[62]=32'h00118903;
    data[63]=32'h00112020;
    data[64]=32'h20020022;
    data[65]=32'h0000000c;
    data[66]=32'h00118903;
    data[67]=32'h00112020;
    data[68]=32'h20020022;
    data[69]=32'h0000000c;
    data[70]=32'h00118903;
    data[71]=32'h00112020;
    data[72]=32'h20020022;
    data[73]=32'h0000000c;
    data[74]=32'h20100001;
    data[75]=32'h00109fc0;
    data[76]=32'h00139fc3;
    data[77]=32'h00008021;
    data[78]=32'h2012000c;
    data[79]=32'h24160003;
    data[80]=32'h26100001;
    data[81]=32'h3210000f;
    data[82]=32'h20080008;
    data[83]=32'h20090001;
    data[84]=32'h00139900;
    data[85]=32'h02709825;
    data[86]=32'h00132020;
    data[87]=32'h20020022;
    data[88]=32'h0000000c;
    data[89]=32'h01094022;
    data[90]=32'h1500fff9;
    data[91]=32'h22100001;
    data[92]=32'h2018000f;
    data[93]=32'h02188024;
    data[94]=32'h00108700;
    data[95]=32'h20080008;
    data[96]=32'h20090001;
    data[97]=32'h00139902;
    data[98]=32'h02709825;
    data[99]=32'h00132021;
    data[100]=32'h20020022;
    data[101]=32'h0000000c;
    data[102]=32'h01094022;
    data[103]=32'h1500fff9;
    data[104]=32'h00108702;
    data[105]=32'h02c9b022;
    data[106]=32'h12c00001;
    data[107]=32'h08000050;
    data[108]=32'h00004020;
    data[109]=32'h01084027;
    data[110]=32'h00084400;
    data[111]=32'h3508ffff;
    data[112]=32'h00082021;
    data[113]=32'h20020022;
    data[114]=32'h0000000c;
    data[115]=32'h2010ffff;
    data[116]=32'h20110000;
    data[117]=32'hae300000;
    data[118]=32'h22100001;
    data[118]=32'h22310004;
    data[119]=32'hae300000;
    data[120]=32'h22100001;
    data[121]=32'h22310004;
    data[122]=32'hae300000;
    data[123]=32'h22100001;
    data[124]=32'h22310004;
    data[125]=32'hae300000;
    data[126]=32'h22100001;
    data[127]=32'h22310004;
    data[128]=32'hae300000;
    data[129]=32'h22100001;
    data[130]=32'h22310004;
    data[131]=32'hae300000;
    data[132]=32'h22100001;
    data[133]=32'h22310004;
    data[134]=32'hae300000;
    data[135]=32'h22100001;
    data[136]=32'h22310004;
    data[137]=32'hae300000;
    data[138]=32'h22100001;
    data[139]=32'h22310004;
    data[140]=32'hae300000;
    data[141]=32'h22100001;
    data[142]=32'h22310004;
    data[143]=32'hae300000;
    data[144]=32'h22100001;
    data[145]=32'h22310004;
    data[146]=32'hae300000;
    data[147]=32'h22100001;
    data[148]=32'h22310004;
    data[149]=32'hae300000;
    data[150]=32'h22100001;
    data[151]=32'h22310004;
    data[152]=32'hae300000;
    data[153]=32'h22100001;
    data[154]=32'h22310004;
    data[155]=32'hae300000;
    data[156]=32'h22100001;
    data[157]=32'h22310004;
    data[158]=32'hae300000;
    data[159]=32'h22100001;
    data[160]=32'h22310004;
    data[161]=32'hae300000;
    data[162]=32'h22100001;
    data[163]=32'h22310004;
    data[164]=32'h22100001;
    data[165]=32'h00008020;
    data[166]=32'h2011003c;
    data[167]=32'h8e130000;
    data[168]=32'h8e340000;
    data[169]=32'h0274402a;
    data[170]=32'h11000002;
    data[171]=32'hae330000;
    data[172]=32'hae140000;
    data[173]=32'h2231fffc;
    data[174]=32'h1611fff8;
    data[175]=32'h00102020;
    data[176]=32'h20020022;
    data[177]=32'h0000000c;
    data[178]=32'h22100004;
    data[179]=32'h2011003c;
    data[180]=32'h1611fff2;
    data[181]=32'h2002000a;
    data[182]=32'h0000000c;
    data[183]=32'h20100000;
    data[184]=32'h22100001;
    data[185]=32'h00102020;
    data[186]=32'h20020022;
    data[187]=32'h0000000c;
    data[188]=32'h22100002;
    data[189]=32'h00102020;
    data[190]=32'h20020022;
    data[191]=32'h0000000c;
    data[192]=32'h22100003;
    data[193]=32'h00102020;
    data[194]=32'h20020022;
    data[195]=32'h0000000c;
    data[196]=32'h22100004;
    data[197]=32'h00102020;
    data[198]=32'h20020022;
    data[199]=32'h0000000c;
    data[200]=32'h22100005;
    data[201]=32'h00102020;
    data[202]=32'h20020022;
    data[203]=32'h0000000c;
    data[204]=32'h22100006;
    data[205]=32'h00102020;
    data[206]=32'h20020022;
    data[207]=32'h0000000c;
    data[208]=32'h22100007;
    data[209]=32'h00102020;
    data[210]=32'h20020022;
    data[211]=32'h0000000c;
    data[212]=32'h22100008;
    data[213]=32'h00102020;
    data[214]=32'h20020022;
    data[215]=32'h20020022;
    data[216]=32'h0000000c;
    data[217]=32'h03e00008;
    end
    always @(address)
    begin
    dataout=data[address];
    end
endmodule
